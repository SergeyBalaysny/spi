library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package parameters is

	constant c_LEN: natural := 127;

end package ; -- parameters_p 
